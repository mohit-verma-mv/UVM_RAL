interface top_if();
  
  logic clk;
  logic rst;
  logic wr;
  logic addr;
  logic [7:0] din;
  logic [7:0] dout;
  
endinterface